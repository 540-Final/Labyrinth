`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/07/2014 05:37:46 PM
// Design Name: 
// Module Name: ball_collision_test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ball_collision_test(
    
   Ball ball
(
	map_value,	
	.clk,
	.reset,	
	.movement,	
	.y_out,
	.x_out,
	
	.vid_row,		// video logic row address
	.vid_col,		// video logic column address
	.vid_pixel_out	// pixel (location) value
);
    
    );
endmodule
